* /home/kanish/eSim-2.3/library/SubcircuitLibrary/cmos_switch_sub/cmos_switch_sub.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Wed Nov 30 22:07:16 2022

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
SC1  A1 Net-_SC1-Pad2_ Vdd Vdd sky130_fd_pr__pfet_01v8_hvt		
SC2  A1 Net-_SC1-Pad2_ gnd gnd sky130_fd_pr__nfet_01v8		
SC5  A2 A1 Vdd Vdd sky130_fd_pr__pfet_01v8_hvt		
SC6  A2 A1 gnd gnd sky130_fd_pr__nfet_01v8		
SC3  Net-_SC3-Pad1_ A1 Net-_SC3-Pad3_ Vdd sky130_fd_pr__pfet_01v8_hvt		
SC8  Net-_SC4-Pad3_ A2 Net-_SC3-Pad1_ Vdd sky130_fd_pr__pfet_01v8_hvt		
SC4  Net-_SC3-Pad1_ A1 Net-_SC4-Pad3_ gnd sky130_fd_pr__nfet_01v8		
SC7  Net-_SC3-Pad3_ A2 Net-_SC3-Pad1_ gnd sky130_fd_pr__nfet_01v8		
U1  Net-_SC1-Pad2_ Net-_SC4-Pad3_ Net-_SC3-Pad3_ Net-_SC3-Pad1_ Vdd gnd PORT		

.end
